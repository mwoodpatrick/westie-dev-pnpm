## @param wordpressUsername WordPress username
##
wordpressUsername: "wp-admin"
wordpressPassword: "wp4MrktOuse1982"
wordpressPlugins: [ "Google Analytics for WordPress" ]

